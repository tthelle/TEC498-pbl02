module logica_or(A, B, S);
	input [7:0] A, B;
	output [7:0] S;
	
	or or0(S[0], A[0], B[0]);
	or or1(S[1], A[1], B[1]);
	or or2(S[2], A[2], B[2]);
	or or3(S[3], A[3], B[3]);
	or or4(S[4], A[4], B[4]);
	or or5(S[5], A[5], B[5]);
	or or6(S[6], A[6], B[6]);
	or or7(S[7], A[7], B[7]);

endmodule